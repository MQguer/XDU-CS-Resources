library verilog;
use verilog.vl_types.all;
entity fourBitCounterAsync_vlg_vec_tst is
end fourBitCounterAsync_vlg_vec_tst;
