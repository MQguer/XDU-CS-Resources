library verilog;
use verilog.vl_types.all;
entity DffValidation_vlg_vec_tst is
end DffValidation_vlg_vec_tst;
