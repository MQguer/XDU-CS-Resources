library verilog;
use verilog.vl_types.all;
entity One_vlg_check_tst is
    port(
        Ci1             : in     vl_logic;
        S               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end One_vlg_check_tst;
