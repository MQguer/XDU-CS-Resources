library verilog;
use verilog.vl_types.all;
entity clock_vlg_check_tst is
    port(
        pin_name2       : in     vl_logic;
        pin_name3       : in     vl_logic;
        pin_name4       : in     vl_logic;
        pin_name5       : in     vl_logic;
        pin_name6       : in     vl_logic;
        pin_name7       : in     vl_logic;
        pin_name8       : in     vl_logic;
        pin_name10      : in     vl_logic;
        pin_name11      : in     vl_logic;
        pin_name12      : in     vl_logic;
        pin_name13      : in     vl_logic;
        pin_name14      : in     vl_logic;
        pin_name15      : in     vl_logic;
        pin_name16      : in     vl_logic;
        pin_name17      : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end clock_vlg_check_tst;
