library verilog;
use verilog.vl_types.all;
entity Decoder_vlg_vec_tst is
end Decoder_vlg_vec_tst;
