library verilog;
use verilog.vl_types.all;
entity voter_vlg_vec_tst is
end voter_vlg_vec_tst;
