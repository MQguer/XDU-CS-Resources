library verilog;
use verilog.vl_types.all;
entity JKffValidation_vlg_vec_tst is
end JKffValidation_vlg_vec_tst;
