library verilog;
use verilog.vl_types.all;
entity fourB_vlg_check_tst is
    port(
        c4              : in     vl_logic;
        s1              : in     vl_logic;
        s2              : in     vl_logic;
        s3              : in     vl_logic;
        s4              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end fourB_vlg_check_tst;
