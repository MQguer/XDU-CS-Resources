library verilog;
use verilog.vl_types.all;
entity moc_vlg_vec_tst is
end moc_vlg_vec_tst;
