library verilog;
use verilog.vl_types.all;
entity hgh_vlg_sample_tst is
    port(
        in1             : in     vl_logic;
        in2             : in     vl_logic;
        in3             : in     vl_logic;
        in5             : in     vl_logic;
        in6             : in     vl_logic;
        pin_name4       : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end hgh_vlg_sample_tst;
