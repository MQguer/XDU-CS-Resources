library verilog;
use verilog.vl_types.all;
entity fullAdder_vlg_vec_tst is
end fullAdder_vlg_vec_tst;
