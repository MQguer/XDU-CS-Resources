library verilog;
use verilog.vl_types.all;
entity modTen_vlg_vec_tst is
end modTen_vlg_vec_tst;
