library verilog;
use verilog.vl_types.all;
entity fourB_vlg_vec_tst is
end fourB_vlg_vec_tst;
