library verilog;
use verilog.vl_types.all;
entity One_vlg_vec_tst is
end One_vlg_vec_tst;
