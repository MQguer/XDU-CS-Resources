library verilog;
use verilog.vl_types.all;
entity hgh_vlg_vec_tst is
end hgh_vlg_vec_tst;
