library verilog;
use verilog.vl_types.all;
entity fourBitCoparer_vlg_vec_tst is
end fourBitCoparer_vlg_vec_tst;
