library verilog;
use verilog.vl_types.all;
entity fourBitCounterSync_vlg_vec_tst is
end fourBitCounterSync_vlg_vec_tst;
