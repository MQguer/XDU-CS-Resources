library verilog;
use verilog.vl_types.all;
entity fourBitCounterAsync_vlg_sample_tst is
    port(
        CP              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end fourBitCounterAsync_vlg_sample_tst;
