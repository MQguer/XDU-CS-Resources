library verilog;
use verilog.vl_types.all;
entity clock is
    port(
        pin_name2       : out    vl_logic;
        pin_name9       : in     vl_logic;
        pin_name1       : in     vl_logic;
        pin_name3       : out    vl_logic;
        pin_name4       : out    vl_logic;
        pin_name5       : out    vl_logic;
        pin_name6       : out    vl_logic;
        pin_name7       : out    vl_logic;
        pin_name8       : out    vl_logic;
        pin_name11      : out    vl_logic;
        pin_name12      : out    vl_logic;
        pin_name13      : out    vl_logic;
        pin_name14      : out    vl_logic;
        pin_name15      : out    vl_logic;
        pin_name16      : out    vl_logic;
        pin_name10      : out    vl_logic;
        pin_name17      : out    vl_logic
    );
end clock;
