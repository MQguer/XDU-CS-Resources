library verilog;
use verilog.vl_types.all;
entity hgh is
    port(
        o1              : out    vl_logic;
        in1             : in     vl_logic;
        in2             : in     vl_logic;
        pin_name4       : in     vl_logic;
        in3             : in     vl_logic;
        in5             : in     vl_logic;
        in6             : in     vl_logic;
        o2              : out    vl_logic;
        o3              : out    vl_logic;
        o4              : out    vl_logic;
        o5              : out    vl_logic;
        o6              : out    vl_logic;
        o7              : out    vl_logic;
        o8              : out    vl_logic
    );
end hgh;
