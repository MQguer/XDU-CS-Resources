library verilog;
use verilog.vl_types.all;
entity multiplexer_vlg_vec_tst is
end multiplexer_vlg_vec_tst;
