library verilog;
use verilog.vl_types.all;
entity distributor_vlg_vec_tst is
end distributor_vlg_vec_tst;
